module hazard_process(
    
)