module forwarding_unit(
    
)